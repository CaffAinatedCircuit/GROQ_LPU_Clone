* NGSPICE file created from hac_deskew_dut.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt hac_deskew_dut VGND VPWR clk delta_t[0] delta_t[10] delta_t[11] delta_t[12]
+ delta_t[13] delta_t[14] delta_t[15] delta_t[1] delta_t[2] delta_t[3] delta_t[4]
+ delta_t[5] delta_t[6] delta_t[7] delta_t[8] delta_t[9] hac_val[0] hac_val[10] hac_val[11]
+ hac_val[12] hac_val[13] hac_val[14] hac_val[15] hac_val[16] hac_val[17] hac_val[18]
+ hac_val[19] hac_val[1] hac_val[20] hac_val[21] hac_val[22] hac_val[23] hac_val[24]
+ hac_val[25] hac_val[26] hac_val[27] hac_val[28] hac_val[29] hac_val[2] hac_val[30]
+ hac_val[31] hac_val[3] hac_val[4] hac_val[5] hac_val[6] hac_val[7] hac_val[8] hac_val[9]
+ instr_data[0] instr_data[10] instr_data[11] instr_data[12] instr_data[13] instr_data[14]
+ instr_data[15] instr_data[16] instr_data[17] instr_data[18] instr_data[19] instr_data[1]
+ instr_data[20] instr_data[21] instr_data[22] instr_data[23] instr_data[24] instr_data[25]
+ instr_data[26] instr_data[27] instr_data[28] instr_data[29] instr_data[2] instr_data[30]
+ instr_data[31] instr_data[32] instr_data[33] instr_data[34] instr_data[35] instr_data[36]
+ instr_data[37] instr_data[38] instr_data[39] instr_data[3] instr_data[4] instr_data[5]
+ instr_data[6] instr_data[7] instr_data[8] instr_data[9] instr_ready instr_valid
+ link_rx[0] link_rx[10] link_rx[11] link_rx[12] link_rx[13] link_rx[14] link_rx[15]
+ link_rx[16] link_rx[17] link_rx[18] link_rx[19] link_rx[1] link_rx[20] link_rx[21]
+ link_rx[22] link_rx[23] link_rx[24] link_rx[25] link_rx[26] link_rx[27] link_rx[28]
+ link_rx[29] link_rx[2] link_rx[30] link_rx[31] link_rx[32] link_rx[33] link_rx[34]
+ link_rx[35] link_rx[36] link_rx[37] link_rx[38] link_rx[39] link_rx[3] link_rx[40]
+ link_rx[41] link_rx[42] link_rx[43] link_rx[44] link_rx[45] link_rx[46] link_rx[47]
+ link_rx[4] link_rx[5] link_rx[6] link_rx[7] link_rx[8] link_rx[9] link_rx_r link_rx_v
+ link_tx[0] link_tx[10] link_tx[11] link_tx[12] link_tx[13] link_tx[14] link_tx[15]
+ link_tx[16] link_tx[17] link_tx[18] link_tx[19] link_tx[1] link_tx[20] link_tx[21]
+ link_tx[22] link_tx[23] link_tx[24] link_tx[25] link_tx[26] link_tx[27] link_tx[28]
+ link_tx[29] link_tx[2] link_tx[30] link_tx[31] link_tx[32] link_tx[33] link_tx[34]
+ link_tx[35] link_tx[36] link_tx[37] link_tx[38] link_tx[39] link_tx[3] link_tx[40]
+ link_tx[41] link_tx[42] link_tx[43] link_tx[44] link_tx[45] link_tx[46] link_tx[47]
+ link_tx[4] link_tx[5] link_tx[6] link_tx[7] link_tx[8] link_tx[9] link_tx_r link_tx_v
+ phase_status[0] phase_status[1] phase_status[2] phase_status[3] phase_status[4]
+ phase_status[5] phase_status[6] phase_status[7] rst_n sac_val[0] sac_val[10] sac_val[11]
+ sac_val[12] sac_val[13] sac_val[14] sac_val[15] sac_val[16] sac_val[17] sac_val[18]
+ sac_val[19] sac_val[1] sac_val[20] sac_val[21] sac_val[22] sac_val[23] sac_val[24]
+ sac_val[25] sac_val[26] sac_val[27] sac_val[28] sac_val[29] sac_val[2] sac_val[30]
+ sac_val[31] sac_val[3] sac_val[4] sac_val[5] sac_val[6] sac_val[7] sac_val[8] sac_val[9]
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ hac_inst.count\[23\] _0120_ _0584_ _0591_ _0592_ VGND VGND VPWR VPWR _0593_
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0985_ _0169_ _0378_ VGND VGND VPWR VPWR hac_val[11] sky130_fd_sc_hd__xnor2_2
XFILLER_0_172_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1468_ VGND VGND VPWR VPWR _1468_/HI link_tx[44] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_52_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1399_ clknet_3_4__leaf_clk _0032_ rst_n VGND VGND VPWR VPWR hac_inst.count\[8\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0770_ hac_inst.count\[23\] _0104_ _0128_ _0135_ _0129_ VGND VGND VPWR VPWR _0228_
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_141_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1322_ clknet_3_3__leaf_clk _0034_ rst_n VGND VGND VPWR VPWR sac_val[0] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1253_ _0563_ _0573_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_142_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1184_ hac_inst.count\[13\] link_rx[21] VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_79_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0968_ _0372_ _0373_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__and2_2
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0899_ _0333_ _0334_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__nand2_2
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_160_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ hac_inst.count\[31\] hac_offset\[31\] VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0753_ _0209_ _0211_ _0164_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a21o_2
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0684_ hac_offset\[18\] hac_inst.count\[18\] VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_177_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1305_ _0102_ _0621_ _0622_ _0623_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__o31ai_2
X_1236_ link_rx[28] hac_inst.count\[20\] VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__and2b_2
X_1167_ hac_offset\[10\] _0503_ phase_status[0] VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1098_ hac_inst.count\[1\] link_rx[9] VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1021_ sac_val[5] _0396_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__nand2_2
XFILLER_0_163_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0805_ _0242_ _0252_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__and2_2
XFILLER_0_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0736_ _0176_ _0177_ _0178_ _0180_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__or4_2
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0667_ phase_status[0] phase_status[5] phase_status[4] VGND VGND VPWR VPWR _0000_
+ sky130_fd_sc_hd__nor3_2
XFILLER_0_23_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1219_ _0546_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_49_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1004_ _0134_ _0222_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0719_ hac_inst.count\[5\] hac_offset\[5\] VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__and2b_2
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0984_ _0172_ _0208_ _0167_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__o21a_2
XFILLER_0_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1467_ VGND VGND VPWR VPWR _1467_/HI link_tx[43] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_52_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1398_ clknet_3_4__leaf_clk _0031_ rst_n VGND VGND VPWR VPWR hac_inst.count\[7\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_89_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1321_ hac_offset\[31\] _0636_ phase_status[0] VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1252_ _0576_ _0577_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1183_ hac_offset\[12\] _0517_ phase_status[0] VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0967_ hac_inst.count\[30\] _0371_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__nand2_2
XFILLER_0_104_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0898_ _0330_ _0332_ _0333_ _0329_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_93_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0821_ _0263_ _0269_ _0270_ _0267_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o31a_2
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0752_ _0198_ _0200_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_141_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ hac_inst.count\[19\] hac_offset\[19\] VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__and2b_2
XFILLER_0_177_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1304_ _0102_ hac_offset\[28\] VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__nand2_2
X_1235_ hac_inst.count\[20\] link_rx[28] VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__and2b_2
XFILLER_0_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1166_ _0501_ _0502_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1097_ link_rx[9] hac_inst.count\[1\] VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__and2b_2
XFILLER_0_48_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1020_ _0396_ _0397_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__and2b_2
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0804_ hac_inst.count\[26\] _0113_ _0250_ _0251_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a31o_2
XFILLER_0_181_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0735_ _0180_ _0193_ _0178_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__a21o_2
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0666_ phase_status[5] phase_status[4] VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_126_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1218_ hac_inst.count\[17\] link_rx[25] VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_0_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1149_ _0470_ _0480_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__and2_2
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ _0222_ _0387_ VGND VGND VPWR VPWR hac_val[20] sky130_fd_sc_hd__nor2_2
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0718_ hac_offset\[7\] hac_inst.count\[7\] VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__xor2_2
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0649_ hac_inst.count\[26\] VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ _0171_ _0208_ VGND VGND VPWR VPWR hac_val[10] sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1466_ VGND VGND VPWR VPWR _1466_/HI link_tx[42] sky130_fd_sc_hd__conb_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1397_ clknet_3_4__leaf_clk _0030_ rst_n VGND VGND VPWR VPWR hac_inst.count\[6\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_52_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1320_ _0634_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1251_ link_rx[29] hac_inst.count\[21\] VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2b_2
X_1182_ _0511_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__xor2_2
XFILLER_0_79_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0966_ hac_inst.count\[30\] _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_31_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0897_ _0330_ _0332_ _0329_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a21o_2
XFILLER_0_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1449_ VGND VGND VPWR VPWR _1449_/HI link_tx[25] sky130_fd_sc_hd__conb_1
XFILLER_0_96_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0820_ _0269_ _0271_ VGND VGND VPWR VPWR hac_val[30] sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0751_ _0169_ _0171_ _0203_ _0207_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__and4_2
XFILLER_0_80_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0682_ hac_offset\[19\] hac_inst.count\[19\] VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1303_ _0617_ _0619_ _0620_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__and3_2
X_1234_ hac_offset\[19\] _0561_ phase_status[0] VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1165_ _0491_ _0495_ _0500_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1096_ hac_offset\[0\] phase_status[0] _0440_ _0442_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__o22a_2
XFILLER_0_87_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0949_ _0362_ _0363_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0803_ _0254_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__nand2_2
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0734_ _0191_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0665_ _0125_ _0126_ VGND VGND VPWR VPWR delta_t[0] sky130_fd_sc_hd__nand2_2
XFILLER_0_110_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1217_ link_rx[25] hac_inst.count\[17\] VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_0_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_148_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1148_ _0470_ _0471_ _0480_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__a31o_2
XFILLER_0_48_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1079_ _0429_ _0430_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_157_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1002_ _0139_ _0221_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__and2_2
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0717_ _0174_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__nand2_2
XFILLER_0_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0648_ hac_offset\[24\] VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ _0207_ _0377_ VGND VGND VPWR VPWR hac_val[9] sky130_fd_sc_hd__xor2_2
XFILLER_0_27_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1465_ VGND VGND VPWR VPWR _1465_/HI link_tx[41] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_52_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1396_ clknet_3_1__leaf_clk _0029_ rst_n VGND VGND VPWR VPWR hac_inst.count\[5\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_52_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1250_ hac_inst.count\[21\] link_rx[29] VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__and2b_2
X_1181_ _0489_ _0512_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_78_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0965_ _0370_ _0371_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_31_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0896_ hac_inst.count\[14\] sac_val[14] VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_120_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1448_ VGND VGND VPWR VPWR _1448_/HI link_tx[24] sky130_fd_sc_hd__conb_1
XFILLER_0_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1379_ clknet_3_0__leaf_clk _0091_ rst_n VGND VGND VPWR VPWR hac_offset\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0750_ _0165_ _0166_ _0172_ _0206_ _0168_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__o41a_2
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0681_ hac_offset\[19\] hac_inst.count\[19\] VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__and2b_2
XFILLER_0_40_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1302_ _0617_ _0619_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_32_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1233_ _0559_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__xnor2_2
X_1164_ _0491_ _0495_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__and3_2
XFILLER_0_79_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1095_ phase_status[0] _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0948_ hac_inst.count\[21\] hac_inst.count\[20\] _0355_ _0361_ VGND VGND VPWR VPWR
+ _0363_ sky130_fd_sc_hd__and4_2
XFILLER_0_126_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0879_ sac_val[11] hac_inst.count\[11\] VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__and2b_2
XFILLER_0_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0802_ hac_offset\[28\] hac_inst.count\[28\] VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0733_ hac_offset\[4\] hac_inst.count\[4\] VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0664_ hac_inst.count\[0\] _0101_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__nand2_2
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1216_ link_rx[25] hac_inst.count\[17\] VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_88_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1147_ hac_inst.count\[6\] _0118_ _0478_ _0479_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__a31o_2
XFILLER_0_133_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1078_ sac_val[29] _0427_ sac_val[30] VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1001_ _0385_ _0386_ VGND VGND VPWR VPWR hac_val[19] sky130_fd_sc_hd__nor2_2
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_179_Right_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0716_ hac_inst.count\[6\] hac_offset\[6\] VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_111_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0647_ hac_offset\[4\] VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_176_Left_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0981_ _0202_ _0204_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_15_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1464_ VGND VGND VPWR VPWR _1464_/HI link_tx[40] sky130_fd_sc_hd__conb_1
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1395_ clknet_3_1__leaf_clk _0028_ rst_n VGND VGND VPWR VPWR hac_inst.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_52_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ hac_inst.count\[10\] _0514_ _0513_ _0505_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_182_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0964_ hac_inst.count\[28\] hac_inst.count\[29\] _0369_ VGND VGND VPWR VPWR _0371_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_156_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0895_ _0331_ _0332_ VGND VGND VPWR VPWR delta_t[13] sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1447_ VGND VGND VPWR VPWR _1447_/HI link_tx[23] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_71_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1378_ clknet_3_3__leaf_clk _0090_ rst_n VGND VGND VPWR VPWR hac_offset\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0680_ _0134_ _0137_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__or2_2
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1301_ hac_inst.count\[28\] link_rx[36] VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__xor2_2
X_1232_ _0554_ _0555_ _0552_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_8_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1163_ _0498_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1094_ hac_inst.count\[0\] link_rx[8] VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0947_ hac_inst.count\[20\] _0360_ hac_inst.count\[21\] VGND VGND VPWR VPWR _0362_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0878_ hac_inst.count\[11\] sac_val[11] VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__and2b_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_3_1__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_8
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0801_ hac_offset\[28\] hac_inst.count\[28\] VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__and2b_2
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0732_ _0188_ _0189_ _0181_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a21o_2
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0663_ hac_inst.count\[0\] sac_val[0] VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_40_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1215_ hac_offset\[16\] _0545_ phase_status[0] VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1146_ _0483_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_49_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1077_ sac_val[29] sac_val[30] _0427_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__and3_2
XFILLER_0_48_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ _0143_ _0220_ _0140_ _0142_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0715_ hac_offset\[6\] hac_inst.count\[6\] VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0646_ hac_inst.count\[7\] VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1129_ hac_inst.count\[6\] link_rx[14] VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0980_ _0201_ _0203_ VGND VGND VPWR VPWR hac_val[8] sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1463_ VGND VGND VPWR VPWR _1463_/HI link_tx[39] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1394_ clknet_3_1__leaf_clk _0027_ rst_n VGND VGND VPWR VPWR hac_inst.count\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0963_ hac_inst.count\[28\] _0369_ hac_inst.count\[29\] VGND VGND VPWR VPWR _0370_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0894_ hac_inst.count\[12\] _0116_ _0327_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_70_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1446_ VGND VGND VPWR VPWR _1446_/HI link_tx[22] sky130_fd_sc_hd__conb_1
XFILLER_0_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1377_ clknet_3_3__leaf_clk _0089_ rst_n VGND VGND VPWR VPWR hac_offset\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1300_ _0112_ link_rx[34] _0609_ _0611_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__o311a_2
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1231_ _0557_ _0558_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__nor2_2
X_1162_ link_rx[18] hac_inst.count\[10\] VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__and2b_2
XFILLER_0_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1093_ _0002_ link_rx[8] VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__nor2_2
XFILLER_0_17_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0946_ hac_inst.count\[20\] _0360_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__xor2_2
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0877_ _0315_ _0317_ VGND VGND VPWR VPWR delta_t[10] sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1429_ VGND VGND VPWR VPWR _1429_/HI link_tx[5] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_3_2__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_74_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0800_ hac_inst.count\[28\] hac_offset\[28\] VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_86_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0731_ _0181_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_107_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0662_ _0123_ _0124_ VGND VGND VPWR VPWR hac_val[0] sky130_fd_sc_hd__nand2_2
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1214_ _0541_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__xor2_2
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1145_ _0108_ link_rx[16] VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_49_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ sac_val[29] _0427_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__xor2_2
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0929_ hac_inst.count\[13\] hac_inst.count\[12\] hac_inst.count\[11\] _0349_ VGND
+ VGND VPWR VPWR _0352_ sky130_fd_sc_hd__and4_2
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0714_ hac_inst.count\[9\] hac_offset\[9\] VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__and2b_2
XFILLER_0_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0645_ hac_inst.count\[8\] VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1128_ hac_offset\[5\] _0469_ phase_status[0] VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1059_ sac_val[20] sac_val[21] sac_val[22] _0415_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_81_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1462_ VGND VGND VPWR VPWR _1462_/HI link_tx[38] sky130_fd_sc_hd__conb_1
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1393_ clknet_3_0__leaf_clk _0024_ rst_n VGND VGND VPWR VPWR hac_inst.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_180_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0962_ hac_inst.count\[28\] _0369_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__xor2_2
XFILLER_0_138_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0893_ _0329_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2b_2
XFILLER_0_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1445_ VGND VGND VPWR VPWR _1445_/HI link_tx[21] sky130_fd_sc_hd__conb_1
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1376_ clknet_3_2__leaf_clk _0088_ rst_n VGND VGND VPWR VPWR hac_offset\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1230_ link_rx[27] hac_inst.count\[19\] VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__and2b_2
XFILLER_0_159_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1161_ hac_inst.count\[10\] link_rx[18] VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__and2b_2
XFILLER_0_56_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1092_ phase_status[5] phase_status[4] _0434_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_177_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0945_ _0359_ _0360_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__nor2_2
XFILLER_0_71_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0876_ _0307_ _0316_ _0308_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1428_ VGND VGND VPWR VPWR _1428_/HI link_tx[4] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_147_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1359_ clknet_3_1__leaf_clk _0071_ rst_n VGND VGND VPWR VPWR hac_offset\[2\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_3_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 clknet_3_3__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_6
XFILLER_0_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0730_ hac_inst.count\[3\] hac_offset\[3\] VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_107_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0661_ _0002_ hac_offset\[0\] VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1213_ _0542_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__or2_2
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1144_ _0108_ link_rx[16] VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__and2_2
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1075_ _0427_ _0428_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__and2b_2
XFILLER_0_172_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0928_ hac_inst.count\[12\] _0351_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0859_ _0300_ _0301_ _0298_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_178_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0713_ _0167_ _0170_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0644_ hac_inst.count\[14\] VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1127_ _0467_ _0468_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_101_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1058_ sac_val[21] _0417_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_145_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_154_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_163_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_172_Left_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_181_Left_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1461_ VGND VGND VPWR VPWR _1461_/HI link_tx[37] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_56_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1392_ clknet_3_1__leaf_clk _0013_ rst_n VGND VGND VPWR VPWR hac_inst.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0961_ _0368_ _0369_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__nor2_2
XFILLER_0_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0892_ sac_val[13] hac_inst.count\[13\] VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_70_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1444_ VGND VGND VPWR VPWR _1444_/HI link_tx[20] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_71_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1375_ clknet_3_2__leaf_clk _0087_ rst_n VGND VGND VPWR VPWR hac_offset\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1160_ hac_offset\[9\] _0497_ phase_status[0] VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1091_ phase_status[5] phase_status[4] _0439_ _0435_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__o31a_2
XFILLER_0_56_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0944_ hac_inst.count\[19\] hac_inst.count\[18\] hac_inst.count\[17\] hac_inst.count\[16\]
+ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__and4_2
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ _0304_ _0309_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nor2_2
XFILLER_0_125_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1427_ VGND VGND VPWR VPWR _1427_/HI link_tx[3] sky130_fd_sc_hd__conb_1
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1358_ clknet_3_1__leaf_clk _0070_ rst_n VGND VGND VPWR VPWR hac_offset\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_3_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1289_ hac_inst.count\[27\] link_rx[35] VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__and2b_2
XFILLER_0_78_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload3 clknet_3_4__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0660_ hac_inst.count\[0\] hac_offset\[0\] VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_123_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1212_ link_rx[24] hac_inst.count\[16\] VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__and2b_2
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1143_ hac_offset\[7\] _0482_ phase_status[0] VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1074_ sac_val[26] sac_val[27] _0423_ sac_val[28] VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__a31o_2
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0927_ hac_inst.count\[11\] _0349_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0858_ _0300_ _0301_ VGND VGND VPWR VPWR delta_t[7] sky130_fd_sc_hd__xor2_2
XFILLER_0_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0789_ hac_inst.count\[24\] _0244_ _0239_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a21o_2
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0712_ _0167_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__and2_2
XFILLER_0_53_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0643_ hac_inst.count\[15\] VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1126_ _0458_ _0462_ _0459_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1057_ _0417_ _0418_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__and2_2
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1109_ hac_inst.count\[3\] link_rx[11] VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__and2b_2
XFILLER_0_178_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ VGND VGND VPWR VPWR _1460_/HI link_tx[36] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_56_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1391_ clknet_3_0__leaf_clk _0002_ rst_n VGND VGND VPWR VPWR hac_inst.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0960_ hac_inst.count\[26\] hac_inst.count\[27\] _0367_ VGND VGND VPWR VPWR _0369_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0891_ hac_inst.count\[13\] sac_val[13] VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__and2b_2
XFILLER_0_137_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1443_ VGND VGND VPWR VPWR _1443_/HI link_tx[19] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_71_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1374_ clknet_3_3__leaf_clk _0086_ rst_n VGND VGND VPWR VPWR hac_offset\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_179_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1090_ _0390_ _0391_ _0437_ _0438_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__nor4_2
XFILLER_0_95_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0943_ hac_inst.count\[19\] hac_inst.count\[18\] hac_inst.count\[17\] _0356_ VGND
+ VGND VPWR VPWR _0360_ sky130_fd_sc_hd__and4_2
XFILLER_0_70_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0874_ _0312_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__nand2_2
XFILLER_0_70_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1426_ VGND VGND VPWR VPWR _1426_/HI link_tx[2] sky130_fd_sc_hd__conb_1
XFILLER_0_103_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1357_ clknet_3_0__leaf_clk _0069_ rst_n VGND VGND VPWR VPWR hac_offset\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_173_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1288_ hac_offset\[26\] _0608_ phase_status[0] VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload4 clknet_3_5__leaf_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_12
XFILLER_0_117_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1211_ hac_inst.count\[16\] link_rx[24] VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__and2b_2
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1142_ _0480_ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_49_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1073_ sac_val[26] sac_val[27] sac_val[28] _0423_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__and4_2
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ hac_inst.count\[11\] _0349_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ _0289_ _0294_ _0296_ _0293_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a31o_2
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0788_ hac_offset\[24\] _0238_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__nor2_2
XFILLER_0_141_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1409_ clknet_3_3__leaf_clk _0011_ rst_n VGND VGND VPWR VPWR hac_inst.count\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ hac_inst.count\[10\] hac_offset\[10\] VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0642_ hac_inst.count\[22\] VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1125_ _0464_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_140_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1056_ sac_val[20] _0415_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or2_2
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0909_ hac_inst.count\[3\] _0339_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1108_ _0102_ hac_offset\[2\] _0451_ _0452_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__a22o_2
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1039_ sac_val[11] sac_val[12] _0404_ sac_val[13] VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__a31o_2
XFILLER_0_165_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_86_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ clknet_3_2__leaf_clk _0000_ rst_n VGND VGND VPWR VPWR instr_ready sky130_fd_sc_hd__dfstp_2
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ _0327_ _0328_ VGND VGND VPWR VPWR delta_t[12] sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_97_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1442_ VGND VGND VPWR VPWR _1442_/HI link_tx[18] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_71_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1373_ clknet_3_3__leaf_clk _0085_ rst_n VGND VGND VPWR VPWR hac_offset\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_169_Left_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_178_Left_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0942_ hac_inst.count\[18\] _0358_ hac_inst.count\[19\] VGND VGND VPWR VPWR _0359_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0873_ sac_val[10] hac_inst.count\[10\] VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_153_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1425_ VGND VGND VPWR VPWR _1425_/HI link_tx[1] sky130_fd_sc_hd__conb_1
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1356_ clknet_3_6__leaf_clk _0068_ rst_n VGND VGND VPWR VPWR phase_status[5] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_108_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ _0604_ _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_108_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload5 clknet_3_6__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_8
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ _0539_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__and2_2
X_1141_ hac_inst.count\[6\] _0118_ _0474_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a21bo_2
XTAP_TAPCELL_ROW_88_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1072_ sac_val[27] _0425_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0925_ _0349_ _0350_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0856_ _0298_ _0299_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0787_ _0225_ _0240_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__and2b_2
XFILLER_0_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1408_ clknet_3_3__leaf_clk _0010_ rst_n VGND VGND VPWR VPWR hac_inst.count\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_162_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1339_ clknet_3_7__leaf_clk _0051_ rst_n VGND VGND VPWR VPWR sac_val[17] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0710_ _0165_ _0166_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0641_ hac_offset\[23\] VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_115_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1124_ link_rx[13] hac_inst.count\[5\] VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_140_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1055_ sac_val[20] _0415_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__nand2_2
XFILLER_0_177_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0908_ hac_inst.count\[0\] hac_inst.count\[3\] hac_inst.count\[2\] hac_inst.count\[1\]
+ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__and4_2
XFILLER_0_4_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0839_ sac_val[4] hac_inst.count\[4\] VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__and2b_2
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_123_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1107_ _0447_ _0450_ phase_status[0] VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_132_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1038_ sac_val[11] sac_val[12] sac_val[13] _0404_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__and4_2
XFILLER_0_48_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_150_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1441_ VGND VGND VPWR VPWR _1441_/HI link_tx[17] sky130_fd_sc_hd__conb_1
XFILLER_0_121_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1372_ clknet_3_2__leaf_clk _0084_ rst_n VGND VGND VPWR VPWR hac_offset\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_171_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ hac_inst.count\[18\] _0358_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__xor2_2
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0872_ sac_val[10] hac_inst.count\[10\] VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__and2b_2
XFILLER_0_113_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1424_ VGND VGND VPWR VPWR _1424_/HI link_tx[0] sky130_fd_sc_hd__conb_1
XFILLER_0_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1355_ clknet_3_3__leaf_clk _0067_ rst_n VGND VGND VPWR VPWR phase_status[4] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_147_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ _0601_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_108_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload6 clknet_3_7__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_8
XFILLER_0_172_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1140_ _0477_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nor2_2
X_1071_ _0425_ _0426_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__and2_2
XFILLER_0_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ hac_inst.count\[9\] _0347_ hac_inst.count\[10\] VGND VGND VPWR VPWR _0350_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_154_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0855_ _0109_ sac_val[7] VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__and2_2
XFILLER_0_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0786_ hac_inst.count\[26\] hac_offset\[26\] VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1407_ clknet_3_3__leaf_clk _0009_ rst_n VGND VGND VPWR VPWR hac_inst.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1338_ clknet_3_6__leaf_clk _0050_ rst_n VGND VGND VPWR VPWR sac_val[16] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_162_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1269_ hac_inst.count\[23\] _0120_ _0119_ hac_inst.count\[22\] VGND VGND VPWR VPWR
+ _0592_ sky130_fd_sc_hd__o211a_2
XFILLER_0_127_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0640_ instr_data[17] VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1123_ link_rx[13] hac_inst.count\[5\] VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__and2b_2
XFILLER_0_177_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1054_ _0415_ _0416_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__and2b_2
XFILLER_0_177_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0907_ _0339_ _0340_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0838_ hac_inst.count\[4\] sac_val[4] VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__and2b_2
XFILLER_0_101_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0769_ _0140_ _0142_ _0145_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or4_2
XFILLER_0_101_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1106_ _0447_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1037_ sac_val[12] _0406_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1440_ VGND VGND VPWR VPWR _1440_/HI link_tx[16] sky130_fd_sc_hd__conb_1
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1371_ clknet_3_2__leaf_clk _0083_ rst_n VGND VGND VPWR VPWR hac_offset\[14\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_71_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ _0357_ _0358_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__nor2_2
XFILLER_0_166_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0871_ hac_inst.count\[10\] sac_val[10] VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1423_ VGND VGND VPWR VPWR phase_status[2] _1423_/LO sky130_fd_sc_hd__conb_1
XFILLER_0_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1354_ clknet_3_3__leaf_clk _0066_ rst_n VGND VGND VPWR VPWR phase_status[0] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_147_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1285_ _0599_ _0600_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_108_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_178_Right_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ sac_val[26] _0423_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or2_2
XFILLER_0_88_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0923_ hac_inst.count\[10\] hac_inst.count\[9\] _0347_ VGND VGND VPWR VPWR _0349_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_83_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0854_ _0109_ sac_val[7] VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__nor2_2
XFILLER_0_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0785_ _0240_ _0241_ VGND VGND VPWR VPWR hac_val[25] sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1406_ clknet_3_2__leaf_clk _0008_ rst_n VGND VGND VPWR VPWR hac_inst.count\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_127_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1337_ clknet_3_6__leaf_clk _0049_ rst_n VGND VGND VPWR VPWR sac_val[15] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_162_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1268_ _0581_ _0587_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1199_ _0529_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__or2_2
XFILLER_0_78_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ hac_inst.count\[5\] link_rx[13] VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1053_ sac_val[17] sac_val[18] _0411_ sac_val[19] VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a31o_2
XFILLER_0_177_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0906_ hac_inst.count\[0\] hac_inst.count\[1\] hac_inst.count\[2\] VGND VGND VPWR
+ VPWR _0340_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0837_ _0282_ _0283_ _0280_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__a21o_2
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0768_ _0127_ _0130_ _0136_ _0138_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__nand4_2
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0699_ hac_offset\[13\] hac_inst.count\[13\] VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__and2b_2
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1105_ _0448_ _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__nor2_2
XFILLER_0_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1036_ sac_val[11] _0404_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__xor2_2
XFILLER_0_177_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_73_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_176_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ sac_val[2] sac_val[3] _0393_ sac_val[4] VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__a31o_2
XFILLER_0_147_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ clknet_3_2__leaf_clk _0082_ rst_n VGND VGND VPWR VPWR hac_offset\[13\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_71_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_138_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ _0310_ _0311_ VGND VGND VPWR VPWR delta_t[9] sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1422_ clknet_3_0__leaf_clk _0026_ rst_n VGND VGND VPWR VPWR hac_inst.count\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_1353_ clknet_3_7__leaf_clk _0065_ rst_n VGND VGND VPWR VPWR sac_val[31] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_147_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1284_ hac_inst.count\[24\] _0121_ _0600_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_108_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0999_ _0140_ _0142_ _0143_ _0220_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o211a_2
XFILLER_0_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0922_ hac_inst.count\[9\] _0347_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__xor2_2
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0853_ _0295_ _0297_ VGND VGND VPWR VPWR delta_t[6] sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0784_ hac_inst.count\[24\] _0111_ _0236_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a21o_2
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1405_ clknet_3_2__leaf_clk _0007_ rst_n VGND VGND VPWR VPWR hac_inst.count\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_127_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1336_ clknet_3_6__leaf_clk _0048_ rst_n VGND VGND VPWR VPWR sac_val[14] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_162_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1267_ hac_inst.count\[24\] link_rx[32] VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__xor2_2
X_1198_ link_rx[23] hac_inst.count\[15\] VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__and2b_2
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1121_ hac_offset\[4\] _0463_ phase_status[0] VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1052_ sac_val[17] sac_val[18] sac_val[19] _0411_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and4_2
XFILLER_0_177_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0905_ hac_inst.count\[0\] hac_inst.count\[2\] hac_inst.count\[1\] VGND VGND VPWR
+ VPWR _0339_ sky130_fd_sc_hd__and3_2
XFILLER_0_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0836_ _0282_ _0283_ VGND VGND VPWR VPWR delta_t[3] sky130_fd_sc_hd__xor2_2
XFILLER_0_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0767_ hac_inst.count\[24\] hac_offset\[24\] VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__xor2_2
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0698_ _0153_ _0156_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_181_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1319_ hac_inst.count\[31\] link_rx[39] VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_111_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1104_ link_rx[10] hac_inst.count\[2\] VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__and2b_2
XFILLER_0_75_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1035_ sac_val[11] _0404_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__nand2_2
XFILLER_0_159_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0819_ _0263_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__nor2_2
XFILLER_0_130_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ sac_val[2] sac_val[3] sac_val[4] _0393_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__and4_2
XFILLER_0_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1421_ clknet_3_0__leaf_clk _0025_ rst_n VGND VGND VPWR VPWR hac_inst.count\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_121_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1352_ clknet_3_7__leaf_clk _0064_ rst_n VGND VGND VPWR VPWR sac_val[30] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_147_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1283_ hac_inst.count\[26\] link_rx[34] VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_108_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ _0144_ _0219_ VGND VGND VPWR VPWR hac_val[18] sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0921_ _0347_ _0348_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__nor2_2
XFILLER_0_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0852_ _0289_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__and2_2
XFILLER_0_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0783_ _0238_ _0239_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1404_ clknet_3_2__leaf_clk _0006_ rst_n VGND VGND VPWR VPWR hac_inst.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_166_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1335_ clknet_3_6__leaf_clk _0047_ rst_n VGND VGND VPWR VPWR sac_val[13] sky130_fd_sc_hd__dfrtp_2
X_1266_ hac_offset\[23\] _0589_ phase_status[0] VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_166_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1197_ hac_inst.count\[15\] link_rx[23] VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__and2b_2
XFILLER_0_176_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_175_Left_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1120_ _0460_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1051_ sac_val[18] _0413_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0904_ hac_inst.count\[0\] hac_inst.count\[1\] VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0835_ _0277_ _0279_ _0276_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a21o_2
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0766_ _0127_ _0224_ VGND VGND VPWR VPWR hac_val[23] sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0697_ _0154_ _0155_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_181_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1318_ _0115_ link_rx[38] _0631_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1249_ hac_offset\[20\] _0575_ phase_status[0] VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1103_ hac_inst.count\[2\] link_rx[10] VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__and2b_2
XFILLER_0_89_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1034_ _0404_ _0405_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__and2b_2
XFILLER_0_177_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0818_ _0254_ _0262_ _0264_ _0255_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_114_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0749_ _0202_ _0204_ _0205_ _0173_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__a31o_2
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1017_ sac_val[3] _0395_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_176_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1420_ clknet_3_0__leaf_clk _0023_ rst_n VGND VGND VPWR VPWR hac_inst.count\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1351_ clknet_3_7__leaf_clk _0063_ rst_n VGND VGND VPWR VPWR sac_val[29] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_79_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1282_ hac_offset\[25\] _0603_ phase_status[0] VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0997_ _0149_ _0384_ VGND VGND VPWR VPWR hac_val[17] sky130_fd_sc_hd__xor2_2
XFILLER_0_42_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0920_ hac_inst.count\[7\] _0345_ hac_inst.count\[8\] VGND VGND VPWR VPWR _0348_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_166_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0851_ _0284_ _0287_ _0290_ _0286_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a211o_2
XFILLER_0_24_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0782_ hac_offset\[25\] hac_inst.count\[25\] VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__and2b_2
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1403_ clknet_3_2__leaf_clk _0005_ rst_n VGND VGND VPWR VPWR hac_inst.count\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_166_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1334_ clknet_3_6__leaf_clk _0046_ rst_n VGND VGND VPWR VPWR sac_val[12] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1265_ _0587_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__xor2_2
X_1196_ hac_offset\[14\] _0528_ phase_status[0] VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1050_ _0413_ _0414_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0903_ _0337_ _0338_ VGND VGND VPWR VPWR delta_t[15] sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0834_ _0280_ _0281_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__nor2_2
XFILLER_0_148_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0765_ _0128_ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__nor2_2
XFILLER_0_45_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0696_ hac_offset\[14\] _0107_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__and2_2
XFILLER_0_45_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1317_ phase_status[0] _0631_ _0632_ _0633_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1248_ _0573_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_16_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1179_ link_rx[18] _0504_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__nor2_2
XFILLER_0_116_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1102_ _0441_ _0444_ _0443_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__a21o_2
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1033_ sac_val[8] sac_val[9] _0400_ sac_val[10] VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a31o_2
XFILLER_0_159_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0817_ _0267_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0748_ _0173_ _0205_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__and2b_2
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0679_ _0134_ _0137_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1016_ sac_val[2] _0393_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_176_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1350_ clknet_3_7__leaf_clk _0062_ rst_n VGND VGND VPWR VPWR sac_val[28] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_147_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1281_ _0599_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0996_ _0150_ _0218_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0850_ _0293_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_126_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0781_ hac_inst.count\[25\] hac_offset\[25\] VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__and2b_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1402_ clknet_3_4__leaf_clk _0004_ rst_n VGND VGND VPWR VPWR hac_inst.count\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_166_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1333_ clknet_3_6__leaf_clk _0045_ rst_n VGND VGND VPWR VPWR sac_val[11] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_127_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1264_ _0576_ _0581_ _0583_ link_rx[30] _0105_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__o32a_2
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1195_ _0526_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0979_ _0177_ _0376_ VGND VGND VPWR VPWR hac_val[7] sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0902_ hac_inst.count\[15\] sac_val[15] VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0833_ hac_inst.count\[3\] sac_val[3] VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__and2b_2
XFILLER_0_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0764_ _0133_ _0134_ _0222_ _0132_ _0130_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__o311a_2
XFILLER_0_84_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0695_ hac_offset\[14\] _0107_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__nor2_2
XFILLER_0_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1316_ _0102_ hac_offset\[30\] VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__and2_2
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1247_ _0564_ _0569_ _0571_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__nor3_2
XFILLER_0_155_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1178_ _0484_ _0493_ _0500_ _0506_ _0491_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_67_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1101_ hac_offset\[1\] _0446_ phase_status[0] VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1032_ sac_val[8] sac_val[9] sac_val[10] _0400_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__and4_2
XFILLER_0_49_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0816_ _0115_ hac_offset\[30\] VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__nand2_2
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0747_ hac_offset\[8\] _0108_ _0173_ _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__o31a_2
XFILLER_0_13_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0678_ hac_inst.count\[20\] hac_offset\[20\] VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__and2b_2
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ sac_val[2] _0393_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1280_ _0600_ _0601_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_147_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ _0152_ _0217_ VGND VGND VPWR VPWR hac_val[16] sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0780_ _0236_ _0237_ VGND VGND VPWR VPWR hac_val[24] sky130_fd_sc_hd__nor2_2
XFILLER_0_141_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1401_ clknet_3_4__leaf_clk _0003_ rst_n VGND VGND VPWR VPWR hac_inst.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_126_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1332_ clknet_3_6__leaf_clk _0044_ rst_n VGND VGND VPWR VPWR sac_val[10] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_127_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1263_ hac_inst.count\[23\] link_rx[31] VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__xor2_2
XFILLER_0_39_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1194_ _0518_ _0522_ _0519_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_135_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0978_ _0176_ _0194_ _0174_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_153_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_171_Left_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0901_ _0107_ sac_val[14] _0335_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o21a_2
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_180_Left_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0832_ sac_val[3] hac_inst.count\[3\] VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__and2b_2
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0763_ _0141_ _0143_ _0220_ _0142_ _0139_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0694_ hac_offset\[15\] hac_inst.count\[15\] VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_150_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1315_ _0629_ _0630_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nand2_2
XFILLER_0_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1246_ _0569_ _0571_ _0564_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__o21a_2
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1177_ _0485_ _0496_ _0500_ _0506_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__and4_2
XFILLER_0_91_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1100_ _0441_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1031_ sac_val[9] _0402_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0815_ _0115_ hac_offset\[30\] VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or2_2
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0746_ hac_offset\[9\] hac_inst.count\[9\] VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0677_ _0131_ _0133_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_36_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1229_ hac_inst.count\[19\] link_rx[27] VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__and2b_2
XFILLER_0_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1014_ _0393_ _0394_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ _0183_ _0187_ _0182_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a21o_2
XFILLER_0_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0994_ _0153_ _0383_ VGND VGND VPWR VPWR hac_val[15] sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1400_ clknet_3_4__leaf_clk _0033_ rst_n VGND VGND VPWR VPWR hac_inst.count\[9\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_166_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1331_ clknet_3_5__leaf_clk _0043_ rst_n VGND VGND VPWR VPWR sac_val[9] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_127_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1262_ hac_offset\[22\] _0586_ phase_status[0] VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1193_ _0524_ _0525_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__nand2_2
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0977_ _0176_ _0194_ VGND VGND VPWR VPWR hac_val[6] sky130_fd_sc_hd__xor2_2
XFILLER_0_104_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_182_Right_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0900_ _0335_ _0336_ VGND VGND VPWR VPWR delta_t[14] sky130_fd_sc_hd__and2_2
XFILLER_0_56_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0831_ _0278_ _0279_ VGND VGND VPWR VPWR delta_t[2] sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0762_ _0141_ _0143_ _0220_ _0142_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a31o_2
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0693_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_181_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1314_ _0625_ _0627_ _0629_ _0624_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__a211o_2
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1245_ _0539_ _0540_ _0570_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__a21o_2
XFILLER_0_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1176_ _0509_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__or2_2
XFILLER_0_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1030_ _0402_ _0403_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and2_2
XFILLER_0_88_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0814_ _0265_ _0266_ VGND VGND VPWR VPWR hac_val[29] sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0745_ _0201_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0676_ _0133_ _0134_ _0132_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__o21a_2
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1228_ hac_offset\[18\] _0556_ phase_status[0] VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1159_ _0492_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ sac_val[0] _0392_ sac_val[1] VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0728_ _0123_ _0186_ _0185_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a21o_2
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0659_ link_rx[36] VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0993_ _0156_ _0382_ _0154_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1476_ VGND VGND VPWR VPWR _1476_/HI phase_status[7] sky130_fd_sc_hd__conb_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1330_ clknet_3_6__leaf_clk _0042_ rst_n VGND VGND VPWR VPWR sac_val[8] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_166_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1261_ _0581_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1192_ link_rx[22] hac_inst.count\[14\] VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_79_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0976_ _0196_ _0375_ VGND VGND VPWR VPWR hac_val[5] sky130_fd_sc_hd__xor2_2
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1459_ VGND VGND VPWR VPWR _1459_/HI link_tx[35] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_87_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0830_ _0125_ _0275_ _0274_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__a21o_2
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0761_ _0147_ _0150_ _0218_ _0148_ _0145_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a311o_2
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0692_ hac_offset\[16\] hac_inst.count\[16\] VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_150_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1313_ _0625_ _0627_ _0624_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__a21o_2
X_1244_ _0541_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__nor2_2
XFILLER_0_79_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1175_ link_rx[20] hac_inst.count\[12\] VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__and2b_2
XFILLER_0_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0959_ hac_inst.count\[26\] _0367_ hac_inst.count\[27\] VGND VGND VPWR VPWR _0368_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ _0254_ _0262_ _0255_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__a21o_2
XFILLER_0_181_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0744_ hac_offset\[8\] hac_inst.count\[8\] VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0675_ hac_offset\[20\] hac_inst.count\[20\] VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__and2b_2
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1227_ _0553_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1158_ _0491_ _0494_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and2_2
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1089_ instr_data[29] instr_data[31] instr_data[30] instr_data[28] VGND VGND VPWR
+ VPWR _0438_ sky130_fd_sc_hd__or4b_2
XFILLER_0_47_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Left_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1012_ _0103_ _0390_ _0391_ sac_val[1] sac_val[0] VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__o311a_2
XFILLER_0_88_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_177_Left_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0727_ hac_offset\[1\] hac_inst.count\[1\] VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0658_ link_rx[32] VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_177_Right_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ _0156_ _0382_ VGND VGND VPWR VPWR hac_val[14] sky130_fd_sc_hd__xor2_2
XFILLER_0_172_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1475_ VGND VGND VPWR VPWR _1475_/HI phase_status[6] sky130_fd_sc_hd__conb_1
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1260_ _0576_ _0583_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__nor2_2
XFILLER_0_78_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1191_ hac_inst.count\[14\] link_rx[22] VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0975_ _0110_ hac_inst.count\[4\] _0193_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1458_ VGND VGND VPWR VPWR _1458_/HI link_tx[34] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_87_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1389_ clknet_3_3__leaf_clk _0001_ rst_n VGND VGND VPWR VPWR link_rx_r sky130_fd_sc_hd__dfstp_2
XFILLER_0_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_122_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0760_ _0147_ _0150_ _0218_ _0148_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a31o_2
XFILLER_0_141_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0691_ hac_offset\[16\] hac_inst.count\[16\] VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_150_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1312_ hac_inst.count\[30\] link_rx[38] VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__xor2_2
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1243_ _0544_ _0546_ _0548_ _0566_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__or4_2
X_1174_ hac_inst.count\[12\] link_rx[20] VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__and2b_2
XFILLER_0_79_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0958_ _0112_ _0367_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0889_ _0322_ _0323_ _0326_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__and3_2
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0812_ _0263_ _0264_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__or2_2
XFILLER_0_154_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0743_ hac_offset\[8\] _0108_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__or2_2
XFILLER_0_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0674_ hac_offset\[21\] hac_inst.count\[21\] VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__and2b_2
XFILLER_0_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1226_ _0547_ _0550_ _0548_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__a21o_2
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1157_ _0492_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1088_ _0436_ instr_data[17] instr_valid VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or3b_2
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1011_ _0101_ _0392_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0726_ hac_offset\[1\] hac_inst.count\[1\] VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__and2b_2
XFILLER_0_111_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0657_ link_rx[31] VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1209_ _0535_ _0489_ _0512_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0709_ _0166_ _0167_ _0165_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o21ba_2
XTAP_TAPCELL_ROW_70_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ _0214_ _0379_ _0159_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o21a_2
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1474_ VGND VGND VPWR VPWR _1474_/HI phase_status[3] sky130_fd_sc_hd__conb_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1190_ hac_offset\[13\] _0523_ phase_status[0] VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0974_ _0193_ _0374_ VGND VGND VPWR VPWR hac_val[4] sky130_fd_sc_hd__and2_2
XFILLER_0_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1457_ VGND VGND VPWR VPWR _1457_/HI link_tx[33] sky130_fd_sc_hd__conb_1
X_1388_ clknet_3_0__leaf_clk _0100_ rst_n VGND VGND VPWR VPWR hac_offset\[31\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_87_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0690_ _0146_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__nor2_2
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1311_ hac_offset\[29\] _0628_ phase_status[0] VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux2_1
X_1242_ _0558_ _0567_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ _0102_ hac_offset\[11\] _0507_ _0508_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0957_ _0366_ _0367_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0888_ _0323_ _0326_ _0322_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0811_ hac_inst.count\[29\] _0114_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__and2_2
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0742_ _0198_ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__and2_2
XFILLER_0_141_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0673_ _0131_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1225_ _0553_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1156_ link_rx[17] hac_inst.count\[9\] VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1087_ instr_data[25] instr_data[24] instr_data[27] instr_data[26] VGND VGND VPWR
+ VPWR _0436_ sky130_fd_sc_hd__or4_2
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1010_ _0103_ _0390_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or3_2
XFILLER_0_77_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0725_ _0182_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_38_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0656_ link_rx[30] VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1208_ _0515_ _0535_ _0536_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__o211a_2
X_1139_ link_rx[15] hac_inst.count\[7\] VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_0_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0708_ hac_offset\[10\] hac_inst.count\[10\] VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_111_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0639_ phase_status[0] VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0990_ _0160_ _0381_ VGND VGND VPWR VPWR hac_val[13] sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1473_ VGND VGND VPWR VPWR _1473_/HI phase_status[1] sky130_fd_sc_hd__conb_1
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ _0191_ _0192_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1456_ VGND VGND VPWR VPWR _1456_/HI link_tx[32] sky130_fd_sc_hd__conb_1
X_1387_ clknet_3_0__leaf_clk _0099_ rst_n VGND VGND VPWR VPWR hac_offset\[30\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_87_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1310_ _0626_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_63_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1241_ _0552_ _0557_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nor2_2
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _0499_ _0501_ _0506_ phase_status[0] VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__o31a_2
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ hac_inst.count\[24\] hac_inst.count\[25\] _0365_ VGND VGND VPWR VPWR _0367_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_55_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0887_ _0302_ _0306_ _0325_ _0324_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o31a_2
XFILLER_0_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1439_ VGND VGND VPWR VPWR _1439_/HI link_tx[15] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0810_ hac_inst.count\[29\] _0114_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__nor2_2
XFILLER_0_108_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0741_ hac_offset\[7\] _0109_ _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__o21a_2
XFILLER_0_3_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0672_ hac_inst.count\[21\] hac_offset\[21\] VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__and2b_2
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1224_ hac_inst.count\[18\] link_rx[26] VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1155_ link_rx[17] hac_inst.count\[9\] VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__and2b_2
XFILLER_0_177_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1086_ phase_status[4] _0433_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0939_ hac_inst.count\[17\] hac_inst.count\[16\] _0355_ VGND VGND VPWR VPWR _0358_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0724_ hac_inst.count\[2\] hac_offset\[2\] VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0655_ link_rx[14] VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1207_ _0534_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__or2_2
XFILLER_0_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1138_ hac_inst.count\[7\] link_rx[15] VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_149_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1069_ sac_val[26] _0423_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0707_ hac_inst.count\[11\] hac_offset\[11\] VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__and2b_2
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0638_ sac_val[0] VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1472_ VGND VGND VPWR VPWR _1472_/HI link_tx_v sky130_fd_sc_hd__conb_1
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_101_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0972_ _0188_ _0190_ VGND VGND VPWR VPWR hac_val[3] sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1455_ VGND VGND VPWR VPWR _1455_/HI link_tx[31] sky130_fd_sc_hd__conb_1
X_1386_ clknet_3_0__leaf_clk _0098_ rst_n VGND VGND VPWR VPWR hac_offset\[29\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_87_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1240_ _0547_ _0565_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1171_ _0499_ _0501_ _0506_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0955_ hac_inst.count\[24\] _0365_ hac_inst.count\[25\] VGND VGND VPWR VPWR _0366_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0886_ _0308_ _0309_ _0315_ _0320_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or4b_2
XFILLER_0_42_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ VGND VGND VPWR VPWR _1438_/HI link_tx[14] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1369_ clknet_3_2__leaf_clk _0081_ rst_n VGND VGND VPWR VPWR hac_offset\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0740_ hac_offset\[7\] _0109_ _0174_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a21o_2
XFILLER_0_123_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0671_ _0128_ _0129_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__and2b_2
XFILLER_0_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1223_ link_rx[26] hac_inst.count\[18\] VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_53_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1154_ _0485_ _0489_ _0484_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1085_ phase_status[4] link_tx_r phase_status[5] VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a21o_2
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0938_ hac_inst.count\[17\] _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0869_ _0304_ _0307_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__and2b_2
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0723_ hac_offset\[2\] hac_inst.count\[2\] VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__and2b_2
XFILLER_0_25_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0654_ link_rx[12] VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1206_ _0510_ _0518_ _0519_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1137_ hac_inst.count\[7\] link_rx[15] VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and2b_2
XFILLER_0_149_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1068_ _0423_ _0424_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__and2b_2
XFILLER_0_87_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0706_ hac_offset\[11\] hac_inst.count\[11\] VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__and2b_2
XFILLER_0_41_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0637_ hac_inst.count\[0\] VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_174_Left_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1471_ VGND VGND VPWR VPWR _1471_/HI link_tx[47] sky130_fd_sc_hd__conb_1
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0971_ _0184_ _0187_ VGND VGND VPWR VPWR hac_val[2] sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1454_ VGND VGND VPWR VPWR _1454_/HI link_tx[30] sky130_fd_sc_hd__conb_1
X_1385_ clknet_3_0__leaf_clk _0097_ rst_n VGND VGND VPWR VPWR hac_offset\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1170_ _0504_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__nor2_2
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0954_ hac_inst.count\[24\] _0365_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__xor2_2
XFILLER_0_172_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ _0308_ _0315_ _0316_ _0320_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__or4b_2
XFILLER_0_125_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1437_ VGND VGND VPWR VPWR _1437_/HI link_tx[13] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1368_ clknet_3_4__leaf_clk _0080_ rst_n VGND VGND VPWR VPWR hac_offset\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1299_ _0601_ _0605_ _0615_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__or3_2
XFILLER_0_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0670_ hac_offset\[22\] _0105_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__nand2_2
XFILLER_0_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1222_ hac_offset\[17\] _0551_ phase_status[0] VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1153_ hac_inst.count\[9\] link_rx[17] VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__nand2b_2
X_1084_ phase_status[0] _0433_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0937_ hac_inst.count\[16\] _0355_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0868_ _0308_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_77_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0799_ _0252_ _0253_ VGND VGND VPWR VPWR hac_val[27] sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0722_ hac_offset\[3\] hac_inst.count\[3\] VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__and2b_2
XFILLER_0_53_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0653_ sac_val[12] VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1205_ _0525_ _0529_ _0530_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1136_ _0102_ hac_offset\[6\] _0476_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__a21o_2
XFILLER_0_79_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1067_ sac_val[23] sac_val[24] _0419_ sac_val[25] VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__a31o_2
XFILLER_0_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_87_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0705_ _0157_ _0158_ _0163_ _0159_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__or4b_2
XFILLER_0_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1119_ _0447_ _0450_ _0455_ _0461_ _0454_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a311o_2
XTAP_TAPCELL_ROW_68_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1470_ VGND VGND VPWR VPWR _1470_/HI link_tx[46] sky130_fd_sc_hd__conb_1
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0970_ _0123_ _0186_ VGND VGND VPWR VPWR hac_val[1] sky130_fd_sc_hd__xor2_2
XFILLER_0_138_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1453_ VGND VGND VPWR VPWR _1453_/HI link_tx[29] sky130_fd_sc_hd__conb_1
X_1384_ clknet_3_0__leaf_clk _0096_ rst_n VGND VGND VPWR VPWR hac_offset\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_179_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0953_ _0364_ _0365_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0884_ _0313_ _0319_ _0318_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_70_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1436_ VGND VGND VPWR VPWR _1436_/HI link_tx[12] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1367_ clknet_3_4__leaf_clk _0079_ rst_n VGND VGND VPWR VPWR hac_offset\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ _0572_ _0595_ _0616_ _0594_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__a211o_2
XFILLER_0_78_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_107_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1221_ _0549_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1152_ hac_offset\[8\] _0490_ phase_status[0] VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1083_ link_rx[41] link_rx[40] _0431_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__or4_2
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0936_ hac_inst.count\[16\] hac_inst.count\[15\] hac_inst.count\[14\] _0352_ VGND
+ VGND VPWR VPWR _0356_ sky130_fd_sc_hd__and4_2
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ sac_val[9] hac_inst.count\[9\] VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__and2b_2
XFILLER_0_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0798_ hac_inst.count\[26\] _0113_ _0247_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_141_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1419_ clknet_3_0__leaf_clk _0022_ rst_n VGND VGND VPWR VPWR hac_inst.count\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0721_ _0110_ hac_inst.count\[4\] _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0652_ hac_inst.count\[30\] VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1204_ _0511_ _0521_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__or3_2
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1135_ phase_status[0] _0474_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__and3_2
XFILLER_0_178_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1066_ sac_val[23] sac_val[24] sac_val[25] _0419_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__and4_2
XFILLER_0_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0919_ hac_inst.count\[8\] hac_inst.count\[7\] _0345_ VGND VGND VPWR VPWR _0347_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_71_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0704_ _0161_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__or2_2
XFILLER_0_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1118_ link_rx[10] _0453_ hac_inst.count\[2\] VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1049_ sac_val[17] _0411_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or2_2
XFILLER_0_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_181_Right_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1452_ VGND VGND VPWR VPWR _1452_/HI link_tx[28] sky130_fd_sc_hd__conb_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1383_ clknet_3_0__leaf_clk _0095_ rst_n VGND VGND VPWR VPWR hac_offset\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_161_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0952_ hac_inst.count\[23\] hac_inst.count\[22\] _0363_ VGND VGND VPWR VPWR _0365_
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_60_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0883_ hac_inst.count\[12\] sac_val[12] VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__xor2_2
XFILLER_0_179_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1435_ VGND VGND VPWR VPWR _1435_/HI link_tx[11] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1366_ clknet_3_4__leaf_clk _0078_ rst_n VGND VGND VPWR VPWR hac_offset\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1297_ _0590_ _0602_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__or3_2
XFILLER_0_179_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1220_ _0541_ _0544_ _0543_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1151_ _0485_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__xor2_2
X_1082_ link_rx[43] link_rx[42] link_rx[44] link_rx[45] VGND VGND VPWR VPWR _0432_
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0935_ _0354_ _0355_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0866_ hac_inst.count\[9\] sac_val[9] VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__and2b_2
XFILLER_0_28_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ _0249_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_77_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1418_ clknet_3_0__leaf_clk _0021_ rst_n VGND VGND VPWR VPWR hac_inst.count\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1349_ clknet_3_7__leaf_clk _0061_ rst_n VGND VGND VPWR VPWR sac_val[27] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0720_ hac_offset\[5\] hac_inst.count\[5\] VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__and2b_2
XFILLER_0_107_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0651_ hac_offset\[29\] VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1203_ _0526_ _0531_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__or2_2
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1134_ _0470_ _0473_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__or2_2
XFILLER_0_178_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1065_ sac_val[24] _0421_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0918_ _0109_ _0345_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_151_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0849_ hac_inst.count\[6\] sac_val[6] VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0703_ hac_inst.count\[12\] hac_offset\[12\] VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__and2b_2
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1117_ _0458_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__nand2_2
XFILLER_0_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1048_ sac_val[17] _0411_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_143_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_161_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_170_Left_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1451_ VGND VGND VPWR VPWR _1451_/HI link_tx[27] sky130_fd_sc_hd__conb_1
X_1382_ clknet_3_0__leaf_clk _0094_ rst_n VGND VGND VPWR VPWR hac_offset\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_172_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0951_ hac_inst.count\[22\] _0363_ hac_inst.count\[23\] VGND VGND VPWR VPWR _0364_
+ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_60_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0882_ _0320_ _0321_ VGND VGND VPWR VPWR delta_t[11] sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1434_ VGND VGND VPWR VPWR _1434_/HI link_tx[10] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1365_ clknet_3_1__leaf_clk _0077_ rst_n VGND VGND VPWR VPWR hac_offset\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1296_ _0604_ _0612_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or2_2
XFILLER_0_179_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_176_Right_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ _0462_ _0472_ _0488_ _0487_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__a31o_2
X_1081_ link_rx[46] link_rx[47] link_rx_v VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0934_ hac_inst.count\[15\] hac_inst.count\[14\] _0352_ VGND VGND VPWR VPWR _0355_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0865_ _0302_ _0305_ VGND VGND VPWR VPWR delta_t[8] sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0796_ hac_offset\[27\] hac_inst.count\[27\] VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__and2b_2
XFILLER_0_51_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1417_ clknet_3_0__leaf_clk _0020_ rst_n VGND VGND VPWR VPWR hac_inst.count\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1348_ clknet_3_7__leaf_clk _0060_ rst_n VGND VGND VPWR VPWR sac_val[26] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1279_ hac_inst.count\[25\] link_rx[33] VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__and2b_2
XFILLER_0_74_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0650_ hac_offset\[26\] VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1202_ hac_offset\[15\] _0533_ phase_status[0] VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1133_ _0470_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nand2_2
XFILLER_0_178_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1064_ _0421_ _0422_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__and2_2
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0917_ _0345_ _0346_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__and2b_2
XFILLER_0_71_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0848_ sac_val[6] hac_inst.count\[6\] VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__and2b_2
XFILLER_0_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0779_ _0225_ _0232_ _0234_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__and3_2
XFILLER_0_101_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0702_ hac_offset\[12\] hac_inst.count\[12\] VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__and2b_2
XFILLER_0_123_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1116_ link_rx[12] hac_inst.count\[4\] VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1047_ _0411_ _0412_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__and2b_2
XFILLER_0_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1450_ VGND VGND VPWR VPWR _1450_/HI link_tx[26] sky130_fd_sc_hd__conb_1
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1381_ clknet_3_0__leaf_clk _0093_ rst_n VGND VGND VPWR VPWR hac_offset\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ _0105_ _0363_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_60_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0881_ _0312_ _0317_ _0313_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_137_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1433_ VGND VGND VPWR VPWR _1433_/HI link_tx[9] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1364_ clknet_3_1__leaf_clk _0076_ rst_n VGND VGND VPWR VPWR hac_offset\[7\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_143_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1295_ hac_offset\[27\] _0614_ phase_status[0] VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1080_ sac_val[31] _0429_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__xor2_2
XFILLER_0_99_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0933_ hac_inst.count\[14\] _0352_ hac_inst.count\[15\] VGND VGND VPWR VPWR _0354_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_83_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0864_ _0302_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or2_2
XFILLER_0_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0795_ hac_inst.count\[27\] hac_offset\[27\] VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_70_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1416_ clknet_3_1__leaf_clk _0019_ rst_n VGND VGND VPWR VPWR hac_inst.count\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_177_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1347_ clknet_3_7__leaf_clk _0059_ rst_n VGND VGND VPWR VPWR sac_val[25] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ link_rx[33] hac_inst.count\[25\] VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_27_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1201_ _0531_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1132_ _0462_ _0472_ _0471_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__a21o_2
XFILLER_0_177_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1063_ sac_val[23] _0419_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or2_2
XFILLER_0_76_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ hac_inst.count\[5\] hac_inst.count\[4\] _0341_ hac_inst.count\[6\] VGND VGND
+ VPWR VPWR _0346_ sky130_fd_sc_hd__a31o_2
XFILLER_0_154_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0847_ _0291_ _0292_ VGND VGND VPWR VPWR delta_t[5] sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0778_ _0232_ _0234_ _0225_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_141_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0701_ _0158_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__and2b_2
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1115_ hac_inst.count\[4\] link_rx[12] VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_71_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1046_ sac_val[14] sac_val[15] _0407_ sac_val[16] VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_105_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1029_ sac_val[8] _0400_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1380_ clknet_3_0__leaf_clk _0092_ rst_n VGND VGND VPWR VPWR hac_offset\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ _0318_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__nor2_2
XFILLER_0_82_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1432_ VGND VGND VPWR VPWR _1432_/HI link_tx[8] sky130_fd_sc_hd__conb_1
X_1363_ clknet_3_1__leaf_clk _0075_ rst_n VGND VGND VPWR VPWR hac_offset\[6\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_143_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1294_ _0612_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_158_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Left_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ _0107_ _0352_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0863_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0794_ hac_inst.count\[27\] hac_offset\[27\] VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__and2b_2
XFILLER_0_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1415_ clknet_3_0__leaf_clk _0018_ rst_n VGND VGND VPWR VPWR hac_inst.count\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1346_ clknet_3_7__leaf_clk _0058_ rst_n VGND VGND VPWR VPWR sac_val[24] sky130_fd_sc_hd__dfrtp_2
X_1277_ hac_inst.count\[24\] _0121_ _0597_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_74_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1200_ _0526_ _0527_ _0525_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1131_ _0460_ _0467_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__nor2_2
X_1062_ sac_val[23] _0419_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nand2_2
XFILLER_0_137_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0915_ hac_inst.count\[6\] hac_inst.count\[5\] hac_inst.count\[4\] _0341_ VGND VGND
+ VPWR VPWR _0345_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_116_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0846_ _0284_ _0287_ _0286_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_70_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0777_ _0232_ _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__nand2_2
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1329_ clknet_3_5__leaf_clk _0041_ rst_n VGND VGND VPWR VPWR sac_val[7] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_78_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_104_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_113_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0700_ hac_inst.count\[13\] hac_offset\[13\] VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_128_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1114_ hac_offset\[3\] _0457_ phase_status[0] VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1045_ sac_val[14] sac_val[15] sac_val[16] _0407_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__and4_2
XFILLER_0_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0829_ _0276_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1028_ sac_val[8] _0400_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1431_ VGND VGND VPWR VPWR _1431_/HI link_tx[7] sky130_fd_sc_hd__conb_1
XFILLER_0_121_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1362_ clknet_3_1__leaf_clk _0074_ rst_n VGND VGND VPWR VPWR hac_offset\[5\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_143_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1293_ _0601_ _0604_ _0606_ link_rx[34] _0112_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__o32a_2
XFILLER_0_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0931_ _0352_ _0353_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__and2b_2
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0862_ _0303_ _0304_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__nor2_2
XFILLER_0_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0793_ _0247_ _0248_ VGND VGND VPWR VPWR hac_val[26] sky130_fd_sc_hd__nor2_2
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1414_ clknet_3_0__leaf_clk _0017_ rst_n VGND VGND VPWR VPWR hac_inst.count\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1345_ clknet_3_7__leaf_clk _0057_ rst_n VGND VGND VPWR VPWR sac_val[23] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1276_ hac_offset\[24\] _0598_ phase_status[0] VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1130_ hac_inst.count\[4\] _0117_ _0464_ _0465_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__a31o_2
XFILLER_0_88_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1061_ _0419_ _0420_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__and2b_2
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ hac_inst.count\[5\] _0343_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0845_ _0288_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0776_ _0212_ _0216_ _0227_ _0233_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__a211o_2
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1328_ clknet_3_5__leaf_clk _0040_ rst_n VGND VGND VPWR VPWR sac_val[6] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1259_ _0576_ _0582_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__and2b_2
XFILLER_0_182_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1113_ _0455_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_109_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1044_ sac_val[15] _0409_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_177_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0828_ hac_inst.count\[2\] sac_val[2] VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0759_ _0212_ _0216_ _0152_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a21o_2
XFILLER_0_101_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1027_ _0400_ _0401_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__and2b_2
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1430_ VGND VGND VPWR VPWR _1430_/HI link_tx[6] sky130_fd_sc_hd__conb_1
XFILLER_0_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1361_ clknet_3_1__leaf_clk _0073_ rst_n VGND VGND VPWR VPWR hac_offset\[4\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_143_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ _0609_ _0610_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_160_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0930_ hac_inst.count\[12\] hac_inst.count\[11\] _0349_ hac_inst.count\[13\] VGND
+ VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a31o_2
XFILLER_0_166_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0861_ _0108_ sac_val[8] VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__nor2_2
XFILLER_0_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0792_ _0242_ _0246_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__and2b_2
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1413_ clknet_3_0__leaf_clk _0016_ rst_n VGND VGND VPWR VPWR hac_inst.count\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1344_ clknet_3_6__leaf_clk _0056_ rst_n VGND VGND VPWR VPWR sac_val[22] sky130_fd_sc_hd__dfrtp_2
X_1275_ _0590_ _0596_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1060_ sac_val[20] sac_val[21] _0415_ sac_val[22] VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__a31o_2
XFILLER_0_88_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0913_ _0343_ _0344_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__and2_2
XFILLER_0_83_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0844_ sac_val[5] hac_inst.count\[5\] VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__and2b_2
XFILLER_0_114_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0775_ _0149_ _0151_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__nand2_2
XFILLER_0_105_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1327_ clknet_3_5__leaf_clk _0039_ rst_n VGND VGND VPWR VPWR sac_val[5] sky130_fd_sc_hd__dfrtp_2
X_1258_ _0573_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_127_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1189_ _0521_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1112_ _0447_ _0450_ _0449_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_109_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1043_ _0409_ _0410_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__and2_2
XFILLER_0_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0827_ sac_val[2] hac_inst.count\[2\] VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__and2b_2
XFILLER_0_4_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0758_ _0212_ _0216_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0689_ hac_inst.count\[17\] hac_offset\[17\] VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__and2b_2
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1026_ sac_val[5] sac_val[6] _0396_ sac_val[7] VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__a31o_2
XFILLER_0_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_71_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_182_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1009_ instr_data[21] instr_data[20] instr_data[23] instr_data[22] VGND VGND VPWR
+ VPWR _0391_ sky130_fd_sc_hd__or4_2
XFILLER_0_77_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_118_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ clknet_3_1__leaf_clk _0072_ rst_n VGND VGND VPWR VPWR hac_offset\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1291_ _0610_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_127_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ _0108_ sac_val[8] VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__and2_2
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0791_ _0246_ _0242_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__and2b_2
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1412_ clknet_3_3__leaf_clk _0015_ rst_n VGND VGND VPWR VPWR hac_inst.count\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1343_ clknet_3_6__leaf_clk _0055_ rst_n VGND VGND VPWR VPWR sac_val[21] sky130_fd_sc_hd__dfrtp_2
X_1274_ _0590_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nand2b_2
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0989_ _0161_ _0379_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__nor2_2
XFILLER_0_14_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0912_ hac_inst.count\[4\] _0341_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or2_2
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0843_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0774_ hac_inst.count\[23\] _0104_ _0228_ _0231_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ clknet_3_5__leaf_clk _0038_ rst_n VGND VGND VPWR VPWR sac_val[4] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_179_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1257_ _0563_ _0577_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_127_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1188_ _0511_ _0516_ _0510_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_67_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1111_ _0453_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_109_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1042_ sac_val[14] _0407_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or2_2
XFILLER_0_49_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0826_ _0125_ _0275_ VGND VGND VPWR VPWR delta_t[1] sky130_fd_sc_hd__xor2_2
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0757_ hac_offset\[15\] _0106_ hac_offset\[14\] _0213_ _0215_ VGND VGND VPWR VPWR
+ _0216_ sky130_fd_sc_hd__o221a_2
X_0688_ hac_offset\[17\] hac_inst.count\[17\] VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1309_ hac_inst.count\[28\] _0122_ _0621_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1025_ sac_val[5] sac_val[6] sac_val[7] _0396_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__and4_2
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0809_ _0257_ _0262_ VGND VGND VPWR VPWR hac_val[28] sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_145_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ instr_data[19] instr_data[18] instr_data[16] VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__or3b_2
XFILLER_0_76_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ link_rx[35] hac_inst.count\[27\] VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__and2b_2
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0790_ _0235_ _0243_ _0245_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1411_ clknet_3_3__leaf_clk _0014_ rst_n VGND VGND VPWR VPWR hac_inst.count\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_121_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1342_ clknet_3_6__leaf_clk _0054_ rst_n VGND VGND VPWR VPWR sac_val[20] sky130_fd_sc_hd__dfrtp_2
X_1273_ _0572_ _0595_ _0594_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0988_ _0379_ _0380_ VGND VGND VPWR VPWR hac_val[12] sky130_fd_sc_hd__nor2_2
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_155_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_164_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0911_ hac_inst.count\[4\] _0341_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0842_ hac_inst.count\[5\] sac_val[5] VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__and2b_2
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0773_ _0229_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_180_Right_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_173_Left_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1325_ clknet_3_5__leaf_clk _0037_ rst_n VGND VGND VPWR VPWR sac_val[3] sky130_fd_sc_hd__dfrtp_2
X_1256_ hac_inst.count\[22\] link_rx[30] VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_179_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _0518_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__nand2_2
XFILLER_0_151_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_182_Left_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1110_ link_rx[11] hac_inst.count\[3\] VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_109_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ sac_val[14] _0407_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__nand2_2
XFILLER_0_88_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0825_ hac_inst.count\[1\] sac_val[1] VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0756_ _0157_ _0159_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0687_ hac_offset\[17\] hac_inst.count\[17\] VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and2b_2
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1308_ _0624_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__and2b_2
XFILLER_0_98_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1239_ _0553_ _0559_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_692 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1024_ sac_val[6] _0398_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0808_ _0245_ _0259_ _0261_ _0258_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__a211o_2
XFILLER_0_114_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0739_ _0191_ _0197_ _0195_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ _0223_ _0389_ VGND VGND VPWR VPWR hac_val[22] sky130_fd_sc_hd__nor2_2
XFILLER_0_159_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_692 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1410_ clknet_3_3__leaf_clk _0012_ rst_n VGND VGND VPWR VPWR hac_inst.count\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_131_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1341_ clknet_3_7__leaf_clk _0053_ rst_n VGND VGND VPWR VPWR sac_val[19] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1272_ _0569_ _0593_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__nor2_2
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0987_ _0163_ _0209_ _0211_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__and3_2
XFILLER_0_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0910_ _0341_ _0342_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0841_ _0284_ _0287_ VGND VGND VPWR VPWR delta_t[4] sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_116_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0772_ _0147_ _0150_ _0227_ _0148_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a211o_2
XFILLER_0_144_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1324_ clknet_3_5__leaf_clk _0036_ rst_n VGND VGND VPWR VPWR sac_val[2] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ _0102_ hac_offset\[21\] _0579_ _0580_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_179_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1186_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ _0407_ _0408_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__and2b_2
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0824_ sac_val[1] hac_inst.count\[1\] VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__and2b_2
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0755_ _0158_ _0161_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__or2_2
XFILLER_0_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0686_ _0144_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1307_ link_rx[37] hac_inst.count\[29\] VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1238_ _0548_ _0543_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_168_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1169_ link_rx[19] hac_inst.count\[11\] VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__and2b_2
XFILLER_0_56_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_671 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1023_ _0398_ _0399_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__and2_2
XFILLER_0_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0807_ _0232_ _0234_ _0260_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0738_ _0176_ _0177_ _0192_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0669_ hac_offset\[22\] _0105_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_175_Right_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1006_ _0136_ _0222_ _0130_ _0135_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_92_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1340_ clknet_3_7__leaf_clk _0052_ rst_n VGND VGND VPWR VPWR sac_val[18] sky130_fd_sc_hd__dfrtp_2
X_1271_ _0564_ _0578_ _0591_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ _0209_ _0211_ _0163_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1469_ VGND VGND VPWR VPWR _1469_/HI link_tx[45] sky130_fd_sc_hd__conb_1
XFILLER_0_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ _0285_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0771_ _0141_ _0143_ _0226_ _0142_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_133_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1323_ clknet_3_3__leaf_clk _0035_ rst_n VGND VGND VPWR VPWR sac_val[1] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1254_ _0563_ _0573_ _0578_ phase_status[0] VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_179_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1185_ link_rx[21] hac_inst.count\[13\] VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__and2b_2
XFILLER_0_182_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ hac_inst.count\[31\] _0373_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0823_ _0272_ _0273_ VGND VGND VPWR VPWR hac_val[31] sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0754_ hac_offset\[15\] _0106_ _0107_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a21o_2
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0685_ hac_offset\[18\] hac_inst.count\[18\] VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1306_ hac_inst.count\[29\] link_rx[37] VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__and2b_2
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1237_ _0562_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__nor2_2
X_1168_ hac_inst.count\[11\] link_rx[19] VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and2b_2
XFILLER_0_67_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1099_ _0443_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_177_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1022_ sac_val[5] _0396_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or2_2
XFILLER_0_49_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0806_ _0243_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0737_ _0178_ _0179_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0668_ hac_inst.count\[23\] hac_offset\[23\] VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_179_Left_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1005_ _0136_ _0388_ VGND VGND VPWR VPWR hac_val[21] sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

